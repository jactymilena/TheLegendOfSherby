----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/21/2022 03:01:43 PM
-- Design Name: 
-- Module Name: tile_actor_buffer - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.tuile_package.ALL;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tile_actor_buffer is
    Port ( i_pixel_x    : in STD_LOGIC_VECTOR  (3 downto 0);
           i_pixel_y    : in STD_LOGIC_VECTOR  (3 downto 0);
           i_tile_id    : in STD_LOGIC_VECTOR  (7 downto 0);
           o_color_code : out STD_ULOGIC_VECTOR (3 downto 0));
end tile_actor_buffer;

architecture Behavioral of tile_actor_buffer is

signal test : integer;
signal selected_tile : tableauCouleur;
signal tiles_buffer  : TuilesTableau := (
    (others=> x"0"),
    (   -- LINK DOWN
          TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, x"1", x"1", x"1", TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, x"1", x"1", x"1", x"1", VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , x"1", x"1", x"1", x"1", VERT1_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , x"1", x"1", BEIGE_CC, x"1", VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, TRANS_CC, BEIGE_CC, TRANS_CC
        , x"1", x"1", BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, TRANS_CC
        , x"1", x"1", BRUN_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BEIGE_CC, JAUNE_CC, VERT1_CC, BEIGE_CC, TRANS_CC, TRANS_CC
        , x"1", x"1", BRUN_CC, BRUN_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, x"1", BEIGE_CC, BRUN_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BEIGE_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, BRUN_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, JAUNE_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, VERT1_CC, VERT1_CC, BRUN_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC
    
    ),
    (   -- LINK FRONT
          TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BEIGE_CC, TRANS_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, TRANS_CC, BEIGE_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BEIGE_CC, TRANS_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, TRANS_CC, BEIGE_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, TRANS_CC
        , TRANS_CC, x"1", x"1", x"1", x"1", x"1", BEIGE_CC, BRUN_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC
        , x"1", x"1", JAUNE_CC, JAUNE_CC, x"1", x"1", BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC
        , x"1", JAUNE_CC, x"1", x"1", JAUNE_CC, x"1", x"1", VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, VERT1_CC, VERT1_CC
        , x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", x"1", BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC
        , x"1", x"1", ROUGE_CC, ROUGE_CC, x"1", x"1", x"1", JAUNE_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC
        , x"1", x"1", x"1", x"1", x"1", x"1", x"1", BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, TRANS_CC
        , x"1", JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, x"1", x"1", VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , x"1", x"1", x"1", x"1", x"1", x"1", BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
    ),
    (   -- LINK LEFT
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, BEIGE_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BEIGE_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , BEIGE_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, TRANS_CC, TRANS_CC, VERT1_CC, TRANS_CC, TRANS_CC
        , BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , BEIGE_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC
    ),
 
    (   -- LINK RIGHT
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, BEIGE_CC, VERT1_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, BEIGE_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC
        , TRANS_CC, TRANS_CC, VERT1_CC, TRANS_CC, TRANS_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, BEIGE_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC    
    ),
    
    (   -- LINK TOP
         TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, JAUNE_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BEIGE_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BEIGE_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BEIGE_CC, BEIGE_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, TRANS_CC, BEIGE_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BEIGE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, JAUNE_CC, BEIGE_CC, BEIGE_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BEIGE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, VERT1_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, BEIGE_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1"
        , TRANS_CC, BRUN_CC, BRUN_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, BEIGE_CC, TRANS_CC, TRANS_CC, x"1", x"1"
        , TRANS_CC, BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, JAUNE_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, x"1", x"1", x"1"
        , TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, x"1", x"1", x"1", x"1"
        , TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, x"1", x"1", x"1", x"1", x"1"
        , TRANS_CC, TRANS_CC, VERT1_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, x"1", x"1", x"1", x"1", x"1", TRANS_CC
        , TRANS_CC, BRUN_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BEIGE_CC, x"1", x"1", TRANS_CC, TRANS_CC
        , BRUN_CC, BRUN_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, VERT1_CC, BEIGE_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, VERT1_CC, VERT1_CC, VERT1_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC
    ),
    (   -- SWORD DOWN
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, JAUNE_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
    ),
    (   -- SWORD LEFT
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC
        , GRIS_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, JAUNE_CC, BRUN_CC, VERT1_CC, VERT1_CC
        , TRANS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
    ),
    (   -- SWORD RIGHT
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, TRANS_CC
        , VERT1_CC, VERT1_CC, BRUN_CC, JAUNE_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, BLEU1_CC, GRIS_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, GRIS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
    ),  
    (   -- SWORD UP
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, GRIS_CC, BLEU1_CC, GRIS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, JAUNE_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, VERT1_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
    ),
    (   -- RED HEART
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", x"1", x"1", TRANS_CC, TRANS_CC, TRANS_CC, x"1", x"1", x"1", TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC
        , TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1"
        , TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1"
        , TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1"
        , TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROUGE_CC, ROUGE_CC, ROUGE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROUGE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        
    ),
    (   -- PINK HEART
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", x"1", x"1", TRANS_CC, TRANS_CC, TRANS_CC, x"1", x"1", x"1", TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC
        , TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1"
        , TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1"
        , TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1"
        , TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROSE_CC, ROSE_CC, ROSE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", ROSE_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, x"1", TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
    ),
    (   -- GOOMPA
        TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, BRUN_CC, NOIR_CC, NOIR_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, NOIR_CC, NOIR_CC, BRUN_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BLANC_CC, NOIR_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, NOIR_CC, BLANC_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC
        , TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BLANC_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, BLANC_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BLANC_CC, NOIR_CC, BLANC_CC, BRUN_CC, BRUN_CC, BLANC_CC, NOIR_CC, BLANC_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BLANC_CC, BLANC_CC, BLANC_CC, BRUN_CC, BRUN_CC, BLANC_CC, BLANC_CC, BLANC_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC
        , BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC, BRUN_CC
        , TRANS_CC, BRUN_CC, BRUN_CC, BRUN_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BRUN_CC, BRUN_CC, BRUN_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, NOIR_CC, NOIR_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, NOIR_CC, NOIR_CC, TRANS_CC, TRANS_CC
        , TRANS_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, BEIGE_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, TRANS_CC
        , TRANS_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, TRANS_CC, TRANS_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, TRANS_CC
        , TRANS_CC, TRANS_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, TRANS_CC, TRANS_CC, TRANS_CC, TRANS_CC, NOIR_CC, NOIR_CC, NOIR_CC, NOIR_CC, TRANS_CC, TRANS_CC
    ),
    others =>  (others => x"0")
);
begin
    process(i_pixel_x, i_pixel_y, i_tile_id)
    begin
        selected_tile <= tiles_buffer(to_integer(unsigned(i_tile_id)));
        o_color_code <= selected_tile(to_integer(unsigned(i_pixel_y))* 16 + to_integer(unsigned(i_pixel_x)));
    end process;
    
end Behavioral;
